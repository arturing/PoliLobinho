module unidade_controle(
    input clock,
    input seed,
    input passa,
    
);




parameter INICIAL = 5'd0;
parameter PREPARA_JOGO = 5'd1;


always@(posedge clock) begin
    case()
    endcase
end


endmodule