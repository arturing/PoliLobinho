module fluxo_dados();
endmodule