module unidade_controle();
endmodule